`default_nettype none
`timescale 1ns/1ps

module register_file(clk, //Note - intentionally does not have a reset!
                     wr_ena, wr_addr, wr_data,
                     rd_addr0, rd_data0,
                     rd_addr1, rd_data1);
   // Not parametrizing, these widths are defined by the RISC-V Spec!
   input wire clk;

   // Write channel
   input wire        wr_ena;
   input wire [4:0]  wr_addr;
   input wire [31:0] wr_data;

   // Two read channels
   input wire   [4:0]  rd_addr0, rd_addr1;
   output logic [31:0] rd_data0, rd_data1;

   logic [31:0] x00;
   always_comb x00 = 32'd0; // ties x00 to ground.

   // DON'T DO THIS:
   // logic [31:0] register_file_registers [31:0]
   // CAN'T: because that's a RAM.
   // Works in simulation, fails miserably in synthesis.

   // Hint - use a scripting language if you get tired of copying and pasting
   // the logic 32 times
   // e.g. python: print(",".join(["x%02d"%i for i in range(0,32)]))
   wire [31:0] x01,x02,x03,x04,x05,x06,x07,x08,x09,x10,x11,x12,x13,x14,x15,x16,x17,x18,x19,x20,x21,x22,x23,x24,x25,x26,x27,x28,x29,x30,x31;
endmodule
